library work;
use work.adder_Wbits.all;
